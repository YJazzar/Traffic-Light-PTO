 module NightTime (clk, laneOutput);
   input clk;
   output [7:0] laneOutput;

   
 endmodule